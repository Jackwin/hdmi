module dac (
    input       ref_clk,  // clk is 10 MHz
    input       reset_n,

    output [13:0] dac_data

);

endmodule